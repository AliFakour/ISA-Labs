// systemverlilog header contain the global package
package globals;

	typedef enum logic [3:0] {
		zero, _y, _2y, _3y, _4y, _n4y, _n3y, _n2y, _ny
	} booth_selection_type;

endpackage
